
interface intf();
  
  logic [7:0] a, b;
  logic en;
  logic [3:0] sel;
  logic [15:0] out;
  
endinterface
